module test_of_full_que_shift() 
    red[7:0] back;
    wire[7:0] head;

    reg[1:0] common_selector;

    
endmodule;